module M;
  always_comb a = b;
endmodule
